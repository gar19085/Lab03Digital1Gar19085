module SOP();

//SOP Tabla 01

reg A, B, C;
wire w1, w2, w3, out;

//Compuertas


